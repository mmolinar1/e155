// author: Matthew Molinar
// email: mmolinar@hmc.edu
// date created: 10/25/2025

// key_expansion.sv

/////////////////////////////////////////////
// key_expansion
// generates keys for add_round_key
// NIST FIPS 197 section 5.2
/////////////////////////////////////////////

module key_expansion(input  logic [127:0] state_in,
                     input logic [127:0] key,
                     output logic [127:0] state_out);
    // 

endmodule