// author: Matthew Molinar
// email: mmolinar@hmc.edu
// date created: 10/24/2025

// shift_rows.sv