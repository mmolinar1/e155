// author: Matthew Molinar
// email: mmolinar@hmc.edu
// date created: 09/1/2025